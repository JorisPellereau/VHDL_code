type t_cst_array is array (0 to 63) of std_logic_vector(7 downto 0);
                    constant C_CST_0 : t_cst_array := (
                      0  => x"00",
                      1  => x"3c",
                      2  => x"7e",
                      3  => x"7e",
                      4  => x"7e",
                      5  => x"7e",
                      6  => x"3c",
                      7  => x"00",
                      8  => x"00",
                      9  => x"00",
                      10 => x"02",
                      11 => x"03",
                      12 => x"01",
                      13 => x"03",
                      14 => x"06",
                      15 => x"0c",
                      16 => x"18",
                      17 => x"30",
                      18 => x"60",
                      19 => x"c0",
                      20 => x"80",
                      21 => x"80",
                      22 => x"c0",
                      23 => x"60",
                      24 => x"30",
                      25 => x"18",
                      26 => x"0c",
                      27 => x"06",
                      28 => x"03",
                      29 => x"01",
                      30 => x"03",
                      31 => x"06",
                      32 => x"0c",
                      33 => x"18",
                      34 => x"30",
                      35 => x"60",
                      36 => x"c0",
                      37 => x"80",
                      38 => x"80",
                      39 => x"c0",
                      40 => x"60",
                      41 => x"30",
                      42 => x"18",
                      43 => x"0c",
                      44 => x"06",
                      45 => x"03",
                      46 => x"01",
                      47 => x"03",
                      48 => x"06",
                      49 => x"0c",
                      50 => x"18",
                      51 => x"30",
                      52 => x"60",
                      53 => x"c0",
                      54 => x"80",
                      55 => x"00",
                      56 => x"00",
                      57 => x"3c",
                      58 => x"7e",
                      59 => x"7e",
                      60 => x"7e",
                      61 => x"7e",
                      62 => x"3c",
                      63 => x"00",
                      );
