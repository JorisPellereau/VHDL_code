type t_cst_array is array (0 to 63) of std_logic_vector(7 downto 0);
constant C_CST_0 : t_cst_array := (
  0 => x"ff",
  1 => x"ff",
  2 => x"ff",
  3 => x"ff",
  4 => x"ff",
  5 => x"ff",
  6 => x"ff",
  7 => x"ff",
  8 => x"ff",
  9 => x"ff",
  10 => x"ff",
  11 => x"ff",
  12 => x"ff",
  13 => x"ff",
  14 => x"ff",
  15 => x"ff",
  16 => x"ff",
  17 => x"ff",
  18 => x"ff",
  19 => x"ff",
  20 => x"ff",
  21 => x"ff",
  22 => x"ff",
  23 => x"ff",
  24 => x"ff",
  25 => x"ff",
  26 => x"ff",
  27 => x"ff",
  28 => x"ff",
  29 => x"ff",
  30 => x"ff",
  31 => x"ff",
  32 => x"ff",
  33 => x"ff",
  34 => x"ff",
  35 => x"ff",
  36 => x"ff",
  37 => x"ff",
  38 => x"ff",
  39 => x"ff",
  40 => x"ff",
  41 => x"ff",
  42 => x"ff",
  43 => x"ff",
  44 => x"ff",
  45 => x"ff",
  46 => x"ff",
  47 => x"ff",
  48 => x"ff",
  49 => x"ff",
  50 => x"ff",
  51 => x"ff",
  52 => x"ff",
  53 => x"ff",
  54 => x"ff",
  55 => x"ff",
  56 => x"ff",
  57 => x"ff",
  58 => x"ff",
  59 => x"ff",
  60 => x"ff",
  61 => x"ff",
  62 => x"fe",
  63 => x"ff"
);