type t_cst_array is array (0 to 63) of std_logic_vector(7 downto 0);
constant C_CST_0 : t_cst_array := (
  0 => x"ff",
  1 => x"c3",
  2 => x"81",
  3 => x"81",
  4 => x"81",
  5 => x"81",
  6 => x"c3",
  7 => x"ff",
  8 => x"ff",
  9 => x"ff",
  10 => x"fd",
  11 => x"fc",
  12 => x"fe",
  13 => x"fc",
  14 => x"f9",
  15 => x"f3",
  16 => x"e7",
  17 => x"cf",
  18 => x"9f",
  19 => x"3f",
  20 => x"7f",
  21 => x"7f",
  22 => x"3f",
  23 => x"9f",
  24 => x"cf",
  25 => x"e7",
  26 => x"f3",
  27 => x"f9",
  28 => x"fc",
  29 => x"fe",
  30 => x"fc",
  31 => x"f9",
  32 => x"f3",
  33 => x"e7",
  34 => x"cf",
  35 => x"9f",
  36 => x"3f",
  37 => x"7f",
  38 => x"7f",
  39 => x"3f",
  40 => x"9f",
  41 => x"cf",
  42 => x"e7",
  43 => x"f3",
  44 => x"f9",
  45 => x"fc",
  46 => x"fe",
  47 => x"fc",
  48 => x"f9",
  49 => x"f3",
  50 => x"e7",
  51 => x"cf",
  52 => x"9f",
  53 => x"3f",
  54 => x"7f",
  55 => x"ff",
  56 => x"ff",
  57 => x"c3",
  58 => x"81",
  59 => x"81",
  60 => x"81",
  61 => x"81",
  62 => x"c3",
  63 => x"ff",
);