type t_cst_array is array (0 to 3) of std_logic_vector(7 downto 0);

                    constant C_CST_0 : t_cst_array := (

                      0 => x"EE",
                      1 => x"FF"

                      );
