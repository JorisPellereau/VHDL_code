-------------------------------------------------------------------------------
-- Title      : PWM command
-- Project    : 
-------------------------------------------------------------------------------
-- File       : pwm.vhd
-- Author     :   <JorisPC@JORISP>
-- Company    : 
-- Created    : 2019-06-19
-- Last update: 2019-06-19
-- Platform   : 
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description: This is a simple PWM command
-------------------------------------------------------------------------------
-- Copyright (c) 2019 
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2019-06-19  1.0      JorisPC	Created
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

