-------------------------------------------------------------------------------
-- Title      : Test of the I2C EEPROM Controller
-- Project    : 
-------------------------------------------------------------------------------
-- File       : test_master_i2c_24lc02b.vhd
-- Author     :   <JorisPC@JORISP>
-- Company    : 
-- Created    : 2019-06-25
-- Last update: 2019-06-25
-- Platform   : 
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description: This is a test
-------------------------------------------------------------------------------
-- Copyright (c) 2019 
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2019-06-25  1.0      JorisPC Created
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

library lib_i2c;
use lib_i2c.pkg_i2c.all;

entity test_master_i2c_24c02b is

end entity test_master_i2c_24c02b;

architecture arch_test_master_i2c_24lc02b of test_master_i2c_24c02b is

begin  -- architecture arch_test_master_i2c_24lc02b



end architecture arch_test_master_i2c_24lc02b;

