-------------------------------------------------------------------------------
-- Title      : ADV7123 interface
-- Project    : 
-------------------------------------------------------------------------------
-- File       : adv7123.vhd
-- Author     : Linux-JP  <linux-jp@linuxjp>
-- Company    : 
-- Created    : 2023-08-02
-- Last update: 2023-08-03
-- Platform   : 
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description: 
-------------------------------------------------------------------------------
-- Copyright (c) 2023 
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2023-08-02  1.0      linux-jp	Created
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

entity adv7123 is
  
  port (
    clk   : in std_logic;               -- Clock in
    rst_n : in std_logic);              -- Asynchronous Reset

end entity adv7123;

architecture rtl of adv7123 is

begin  -- architecture rtl

  

end architecture rtl;
