-------------------------------------------------------------------------------
-- Title      : Pseudo Random Binary Sequence Package
-- Project    : 
-------------------------------------------------------------------------------
-- File       : pkg_prbs.vhd
-- Author     :   <JorisPC@JORISP>
-- Company    : 
-- Created    : 2019-06-03
-- Last update: 2019-06-03
-- Platform   : 
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description: This is the package of the PRBS
-------------------------------------------------------------------------------
-- Copyright (c) 2019 
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2019-06-03  1.0      JorisPC Created
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

library lib_prbs;
use lib_prbs.pkg_prbs.all;

package pkg_prbs is

  type int_array is array(0 to 3) of integer range 0 to 32;
  type prbs_features is record
    prbs_alias   : string(1 to 6);
    lfsr_size    : integer range 2 to 32;
    fbk_number   : integer range 2 to 4;
    fbk_position : int_array;
  end record;

  type prbs_type is array(2 to 32) of prbs_features;


  constant prbs_cst : prbs_type := (
    2  => ("PRBS02", 2, 2, (0, 1, 0, 0)),  -- x^2 + X + 1
    3  => ("PRBS03", 3, 2, (0, 1, 0, 0)),  -- X^3 + X + 1                        
    4  => ("PRBS04", 4, 2, (0, 1, 0, 0)),  -- X^4 + X^3 + 1
    5  => ("PRBS05", 5, 2, (0, 2, 0, 0)),  -- X^5 + X^3 + 1
    6  => ("PRBS06", 6, 2, (0, 1, 0, 0)),  -- X^6 + X^5 + 1
    7  => ("PRBS07", 7, 2, (0, 1, 0, 0)),  -- X^7 + X^6 + 1
    8  => ("PRBS08", 8, 4, (0, 2, 3, 4)),  -- X^8 + X^6 + X^5 + X^4 + 1
    9  => ("PRBS09", 9, 2, (0, 4, 0, 0)),  -- X^9 + X^5 + 1
    10 => ("PRBS10", 10, 2, (0, 3, 0, 0)),     -- X^10 + X^7 + 1
    11 => ("PRBS11", 11, 2, (0, 2, 0, 0)),     -- X^11 + X^9 + 1
    12 => ("PRBS12", 12, 4, (0, 6, 8, 11)),    -- X^12 + X^6 + X^4 + X + 1
    13 => ("PRBS13", 13, 4, (0, 9, 10, 12)),   -- X^13 + X^4 + X^3 + X + 1
    14 => ("PRBS14", 14, 4, (0, 9, 11, 13)),   -- X^14 + X^5 + X^3 + X + 1
    15 => ("PRBS15", 15, 2, (0, 1, 0, 0)),     -- X^15 + X^14 + 1
    16 => ("PRBS16", 16, 4, (0, 1, 3, 12)),    -- X^16 + X^15 + X^13 + X^4 + 1
    17 => ("PRBS17", 17, 2, (0, 3, 0, 0)),     -- X^17 + X^14 + 1
    18 => ("PRBS18", 18, 2, (0, 7, 0, 0)),     -- X^18 + X^11 + 1
    19 => ("PRBS19", 19, 4, (0, 13, 17, 18)),  -- X^19 + X^6 + X^2 + X + 1
    20 => ("PRBS20", 20, 2, (0, 3, 0, 0)),     -- X^20 + X^17 + 1
    21 => ("PRBS21", 21, 2, (0, 2, 0, 0)),     -- X^21 + X^19 + 1
    22 => ("PRBS22", 22, 2, (0, 1, 0, 0)),     -- X^22 + X^21 + 1
    23 => ("PRBS23", 23, 2, (0, 5, 0, 0)),     -- X^23 + X^18 + 1
    24 => ("PRBS24", 24, 4, (0, 1, 2, 7)),     -- X^24 + X^23 + X^22 + X^17 + 1
    25 => ("PRBS25", 25, 2, (0, 3, 0, 0)),     -- X^25 + X^22 + 1
    26 => ("PRBS26", 26, 4, (0, 20, 24, 25)),  -- X^26 + X^6 + X^2 + X + 1
    27 => ("PRBS27", 27, 4, (0, 22, 25, 26)),  -- X^27 + X^5 + X^2 + X + 1
    28 => ("PRBS28", 28, 2, (0, 3, 0, 0)),     -- X^28 + X^25 + 1
    29 => ("PRBS29", 29, 2, (0, 2, 0, 0)),     -- X^29 + X^27 + 1
    30 => ("PRBS30", 30, 4, (0, 24, 26, 29)),  -- X^30 + X^6 + X^4 + X + 1
    31 => ("PRBS31", 31, 2, (0, 3, 0, 0)),     -- X^31 + X^28 + 1
    32 => ("PRBS32", 32, 4, (0, 10, 30, 31))   -- X^32 + x^22 + X + X + 1
    );

  component prbs is
    generic(
      prbs_i : integer range 2 to 32 := 3  -- PRBS index 2 => 32
      );
    port(
      -- == INPUTS ==
      lfsr_preload : in  std_logic_vector(prbs_cst(prbs_i).lfsr_size - 1 downto 0);  -- Preload of the LFSR
      clk          : in  std_logic;     -- Clock
      rst_n        : in  std_logic;     -- Asynchron RESET
      start        : in  std_logic;     -- Start the sequence
      -- == OUTPUTS ==
      lfsr         : out std_logic_vector(prbs_cst(prbs_i).lfsr_size - 1 downto 0);  -- LFSR output
      d_out        : out std_logic      -- Serial output
      );
  end component;


end pkg_prbs;

--constant prbs_cst : prbs_type := (
--      2       => ("PRBS02", 2 , 2 , (2 , 1 , 0 , 0)),                                         --
--      3       => ("PRBS03", 3 , 2 , (3 , 2 , 0 , 0)),                                                         
--      4       => ("PRBS04", 4 , 2 , (4 , 3 , 0 , 0)),
--      5       => ("PRBS05", 5 , 2 , (5 , 3 , 0 , 0)),
--      6       => ("PRBS06", 6 , 2 , (6 , 5 , 0 , 0)),
--      7       => ("PRBS07", 7 , 2 , (7 , 6 , 0 , 0)),
--      8       => ("PRBS08", 8 , 4 , (8 , 6 , 5 , 4)),
--      9       => ("PRBS09", 9 , 2 , (9 , 5 , 0 , 0)),
--      10      => ("PRBS10", 11 , 2 , (10 , 7 , 0 , 0)),
--      11      => ("PRBS11", 10 , 2 , (11 , 9 , 0 , 0)),
--      12      => ("PRBS12", 12 , 4 , (12 , 6 , 4 , 1)),
--      13      => ("PRBS13", 13 , 4 , (13 , 4 , 3 , 1)),
--      14      => ("PRBS14", 14 , 4 , (14 , 5 , 3 , 1)),
--      15      => ("PRBS15", 15 , 2 , (15 , 14 , 0 , 0)),
--      16      => ("PRBS16", 16 , 4 , (16 , 15 , 13 , 4)),
--      17      => ("PRBS17", 17 , 2 , (17 , 14 , 0 , 0)),
--      18      => ("PRBS18", 18 , 2 , (18 , 11 , 0 , 0)),
--      19      => ("PRBS19", 19 , 4 , (19 , 6 , 2 , 1)),
--      20      => ("PRBS20", 20 , 2 , (20 , 17 , 0 , 0)),
--      21      => ("PRBS21", 21 , 2 , (21 , 19 , 0 , 0)),
--      22      => ("PRBS22", 22 , 2 , (22 , 21 , 0 , 0)),
--      23      => ("PRBS23", 23 , 2 , (23 , 18 , 0 , 0)),
--      24      => ("PRBS24", 24 , 4 , (24 , 23 , 22 , 17)),
--      25      => ("PRBS25", 25 , 2 , (25 , 22 , 0 , 0)),
--      26      => ("PRBS26", 26 , 4 , (26 , 6 , 2 , 1)),
--      27      => ("PRBS27", 27 , 4 , (27 , 5 , 2 , 1)),
--      28      => ("PRBS28", 28 , 2 , (28 , 25 , 0 , 0)),
--      29      => ("PRBS29", 29 , 2 , (29 , 27 , 0 , 0)),
--      30      => ("PRBS30", 30 , 4 , (30 , 6 , 4 ,  1)),
--      31      => ("PRBS31", 31 , 2 , (31 , 28 , 0 , 0)),
--      32      => ("PRBS32", 32 , 4 , (32 , 22 , 2 , 1))
--);

